// lms_dsp_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module lms_dsp_tb (
	);

	wire         lms_dsp_inst_clk_bfm_clk_clk;                     // lms_dsp_inst_clk_bfm:clk -> [lms_dsp_inst:clk_clk, lms_dsp_inst_fifo_in_bfm:clk, lms_dsp_inst_fifo_out_bfm:clk, lms_dsp_inst_ppd_bfm:clk, lms_dsp_inst_reset_bfm:clk]
	wire   [0:0] lms_dsp_inst_fifo_in_bfm_conduit_wrreq;           // lms_dsp_inst_fifo_in_bfm:sig_wrreq -> lms_dsp_inst:fifo_in_wrreq
	wire  [47:0] lms_dsp_inst_fifo_in_bfm_conduit_wdata;           // lms_dsp_inst_fifo_in_bfm:sig_wdata -> lms_dsp_inst:fifo_in_wdata
	wire         lms_dsp_inst_fifo_out_wrreq;                      // lms_dsp_inst:fifo_out_wrreq -> lms_dsp_inst_fifo_out_bfm:sig_wrreq
	wire  [47:0] lms_dsp_inst_fifo_out_wrdata;                     // lms_dsp_inst:fifo_out_wrdata -> lms_dsp_inst_fifo_out_bfm:sig_wrdata
	wire   [0:0] lms_dsp_inst_ppd_bfm_conduit_cfg_clear_rs;        // lms_dsp_inst_ppd_bfm:sig_cfg_clear_rs -> lms_dsp_inst:ppd_cfg_clear_rs
	wire  [31:0] lms_dsp_inst_ppd_debug_count;                     // lms_dsp_inst:ppd_debug_count -> lms_dsp_inst_ppd_bfm:sig_debug_count
	wire   [0:0] lms_dsp_inst_ppd_bfm_conduit_cfg_enable;          // lms_dsp_inst_ppd_bfm:sig_cfg_enable -> lms_dsp_inst:ppd_cfg_enable
	wire  [31:0] lms_dsp_inst_ppd_debug_long_sum;                  // lms_dsp_inst:ppd_debug_long_sum -> lms_dsp_inst_ppd_bfm:sig_debug_long_sum
	wire   [7:0] lms_dsp_inst_ppd_bfm_conduit_cfg_threshold;       // lms_dsp_inst_ppd_bfm:sig_cfg_threshold -> lms_dsp_inst:ppd_cfg_threshold
	wire  [15:0] lms_dsp_inst_ppd_bfm_conduit_cfg_passthrough_len; // lms_dsp_inst_ppd_bfm:sig_cfg_passthrough_len -> lms_dsp_inst:ppd_cfg_passthrough_len
	wire  [31:0] lms_dsp_inst_ppd_debug_short_sum;                 // lms_dsp_inst:ppd_debug_short_sum -> lms_dsp_inst_ppd_bfm:sig_debug_short_sum
	wire         lms_dsp_inst_reset_bfm_reset_reset;               // lms_dsp_inst_reset_bfm:reset -> [lms_dsp_inst:reset_reset_n, lms_dsp_inst_fifo_in_bfm:reset, lms_dsp_inst_fifo_out_bfm:reset, lms_dsp_inst_ppd_bfm:reset]

	lms_dsp lms_dsp_inst (
		.clk_clk                 (lms_dsp_inst_clk_bfm_clk_clk),                     //      clk.clk
		.fifo_in_wdata           (lms_dsp_inst_fifo_in_bfm_conduit_wdata),           //  fifo_in.wdata
		.fifo_in_wrreq           (lms_dsp_inst_fifo_in_bfm_conduit_wrreq),           //         .wrreq
		.fifo_out_wrdata         (lms_dsp_inst_fifo_out_wrdata),                     // fifo_out.wrdata
		.fifo_out_wrreq          (lms_dsp_inst_fifo_out_wrreq),                      //         .wrreq
		.ppd_cfg_passthrough_len (lms_dsp_inst_ppd_bfm_conduit_cfg_passthrough_len), //      ppd.cfg_passthrough_len
		.ppd_cfg_threshold       (lms_dsp_inst_ppd_bfm_conduit_cfg_threshold),       //         .cfg_threshold
		.ppd_cfg_clear_rs        (lms_dsp_inst_ppd_bfm_conduit_cfg_clear_rs),        //         .cfg_clear_rs
		.ppd_cfg_enable          (lms_dsp_inst_ppd_bfm_conduit_cfg_enable),          //         .cfg_enable
		.ppd_debug_count         (lms_dsp_inst_ppd_debug_count),                     //         .debug_count
		.ppd_debug_long_sum      (lms_dsp_inst_ppd_debug_long_sum),                  //         .debug_long_sum
		.ppd_debug_short_sum     (lms_dsp_inst_ppd_debug_short_sum),                 //         .debug_short_sum
		.reset_reset_n           (lms_dsp_inst_reset_bfm_reset_reset)                //    reset.reset_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (125000000),
		.CLOCK_UNIT (1)
	) lms_dsp_inst_clk_bfm (
		.clk (lms_dsp_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm lms_dsp_inst_fifo_in_bfm (
		.clk       (lms_dsp_inst_clk_bfm_clk_clk),           //     clk.clk
		.reset     (~lms_dsp_inst_reset_bfm_reset_reset),    //   reset.reset
		.sig_wdata (lms_dsp_inst_fifo_in_bfm_conduit_wdata), // conduit.wdata
		.sig_wrreq (lms_dsp_inst_fifo_in_bfm_conduit_wrreq)  //        .wrreq
	);

	altera_conduit_bfm_0002 lms_dsp_inst_fifo_out_bfm (
		.clk        (lms_dsp_inst_clk_bfm_clk_clk),        //     clk.clk
		.reset      (~lms_dsp_inst_reset_bfm_reset_reset), //   reset.reset
		.sig_wrdata (lms_dsp_inst_fifo_out_wrdata),        // conduit.wrdata
		.sig_wrreq  (lms_dsp_inst_fifo_out_wrreq)          //        .wrreq
	);

	altera_conduit_bfm_0003 lms_dsp_inst_ppd_bfm (
		.clk                     (lms_dsp_inst_clk_bfm_clk_clk),                     //     clk.clk
		.reset                   (~lms_dsp_inst_reset_bfm_reset_reset),              //   reset.reset
		.sig_cfg_clear_rs        (lms_dsp_inst_ppd_bfm_conduit_cfg_clear_rs),        // conduit.cfg_clear_rs
		.sig_cfg_enable          (lms_dsp_inst_ppd_bfm_conduit_cfg_enable),          //        .cfg_enable
		.sig_cfg_passthrough_len (lms_dsp_inst_ppd_bfm_conduit_cfg_passthrough_len), //        .cfg_passthrough_len
		.sig_cfg_threshold       (lms_dsp_inst_ppd_bfm_conduit_cfg_threshold),       //        .cfg_threshold
		.sig_debug_count         (lms_dsp_inst_ppd_debug_count),                     //        .debug_count
		.sig_debug_long_sum      (lms_dsp_inst_ppd_debug_long_sum),                  //        .debug_long_sum
		.sig_debug_short_sum     (lms_dsp_inst_ppd_debug_short_sum)                  //        .debug_short_sum
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) lms_dsp_inst_reset_bfm (
		.reset (lms_dsp_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (lms_dsp_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
